module main

import tui_console

fn main() {
	tui_console.run()!
}
